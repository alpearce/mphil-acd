#-
# Copyright (c) 2013 Colin Rothwell
# All rights reserved.
#
# This software was developed by Colin Rothwell as part of his final year
# undergraduate project.
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions
# are met:
# 1. Redistributions of source code must retain the above copyright
#    notice, this list of conditions and the following disclaimer.
# 2. Redistributions in binary form must reproduce the above copyright
#    notice, this list of conditions and the following disclaimer in the
#    documentation and/or other materials provided with the distribution.
#
# THIS SOFTWARE IS PROVIDED BY THE AUTHOR AND CONTRIBUTORS ``AS IS'' AND
# ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED.  IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE LIABLE
# FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
# DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
# OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
# HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
# LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
# OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
# SUCH DAMAGE.
#
/*
 * This is currently not working.
 * It needs to be updated to use the server creation stuff, which never quite
 * happened.
 */

import CoProFPServerCreation::*;
import CoProFPMegafunctionSimulation::*;
import CoProFPSimulatedOps::*;
import CoProFPTypes::*;

import MIPS::*;

import List::*;

(* synthesize *)
module mkDiadicMegafunctionWrapperTestBench (Empty);
    List#(MIPSReg) testData =
        cons('h3F800000, //1
        cons('h3F800000,
        cons('h47C35000, //1e5
        cons('h40000000, //2
        cons('h43670000, //231
        cons('h3E2AAA7E, //0.166666
        cons('h41BE8D50, //23.819
        cons('h794F233B, //~6.722e34
        cons('h4C465D40, //5.2e7
        cons('h40000000,
        nil))))))))));
    int testDataCount = fromInteger(length(testData));

    Reg#(Bool) loadingIntoWrapped <- mkReg(False);
    Reg#(int) datumIndex <- mkReg(0);

    SimulatedDiadicMegafunction#(7) addMegafunction 
        <- mkSimulatedDiadicMegafunction(add_fn);
    WrappedMegafunctionALUOpDiad#(7) addWrapper <-
        mkALUOpDiad(addMegafunction.mf);
    CoProFPALUOpDiad wrappedAdd = addWrapper.op;

    rule loadDataIntoRaw (!loadingIntoWrapped);
        let datum = testData[datumIndex];
        rawAdd.load(datum, datum, S, RN);
        if (datumIndex != (testDataCount - 1)) begin
            datumIndex <= datumIndex + 1;
        end
        else begin
            datumIndex <= 0;
            loadingIntoWrapped <= True;
        end
        $display("Loaded Raw result %X", rawAdd.result());
    endrule

    rule loadResultFromRaw;
        $display("Raw result %X", rawAdd.result());
    endrule

    rule loadDataIntoWrapped (loadingIntoWrapped && datumIndex < testDataCount);
        let datum = testData[datumIndex];
        wrappedAdd.load(datum, datum, S, RN);
        datumIndex <= datumIndex + 1;
    endrule

    rule loadResultFromWrapped(loadingIntoWrapped);
        $display("Wrapped result %X", wrappedAdd.result());
    endrule

    rule finish (loadingIntoWrapped && datumIndex == testDataCount);
        $finish();
    endrule
endmodule
