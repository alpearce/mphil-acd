
`define pfcmsizeblg2 17  /* must be at least 16, or change inlined hash function */
`define vdim (1024*64) /* must be a power of two */
`define vfcmsizeblg2 19
`define vdfcmsizeblg2 17
`define PFCMB0SIZE (1<<17)*2 
`define pfcmb2size (1<<(17+2))*2 
`define vdfcmb0size (1<<19)*2
`define vdfcmb2size (1<<(19+2))*2
`define vfcmbsize (1<<19)*2

`define BufElems 8192

`define intsize 32 

